module main

const (
	bread_kinds = [
		'white',
		'wheat',
		'grain',
		'rye',
		'bagel',
		'baguette',
		'pita',
		'ciabatta',
		'focaccia',
	]
)
